module pcie_wr_ctlr (
   input clk ,
   input rst_n  
);

endmodule