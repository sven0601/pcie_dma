module pcie_rd_ctlr (
   input clk ,
   input rst_n  
);

endmodule